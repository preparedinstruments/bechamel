
module vga_sync_test(
    input wire clk_in,
	input wire [8:0] key,
	input wire rpi_vsync,
	input wire rpi_hsync,
	input wire analog_in,
	inout pot_in,
	output [3:0] hdmi_p,
	output [3:0] hdmi_n,
     output reg [3:0] r_out,
     output reg [3:0] b_out,
     output reg [3:0] g_out,
     output wire h_sync,
     output wire v_sync,
     output wire red_led,
	output wire green_led
  );
  
  

//160x120
reg [0:19199] heart =

{
160'b0000000000000000000000000000000000000011111111111111111111111111111111111101111100001111110000011111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000011111111111111111111111111111111111100000111111111111111000011100111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000110000110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000110000011011111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000110000011111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000000001101111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000000111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000001111001111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111,
160'b0000000000000000000000000000000111000001111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000010011001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000001000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000011000000000000000101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000001111110000000011111111001111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000001111111110000011111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000011111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000001111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000001100111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000111111111111111111111111111111101111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000100000111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000111111111111111111111111111111111111111111111101111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000000000111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000110000001111111111111111111111111111111111111111111111110001111111000001111100001111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000001110000001111111111111111111111111111111111111111111111100001111111000001111110001111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000110000000011111111111111111111111111111111111111111111111000000111111100000111111000111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000100000000111111111111111111111111111111111111110111111110000000000000000001111111000000001111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000111111111111111111111111111111111111111110111111111100000000001111111111111110110000111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000000011111101111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000001100000111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000001100011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000001100011111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000110011111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000001110111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000011110011111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000111111011111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1000111011111111111111111111111111111111111111111111111111111110001111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1100100000001111111111110111111111111111111111111110111111111100001111111111110000111011111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1100000000000111111110011111111111111111111111111100111111111100001111111111110000010001111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1000000000000111111100011111111111111111111111111000111111111000000111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1000000000000111111100111111111111111111111111111100111111111100010111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0000000000001111111111111111111111111111111111111111111111111111110111111111000110000100111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0111000000000111111111111111111111111111111111110110011111111111111111100010001111111110011111111111111111111111111111111111111111111111111111111111111111111111,
160'b0111100000000001011111111111111111111111111111111110011111111111101111000000001111111110001111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111110000000000011111111111111111111111111111111111011111111111100110000000000110000000011111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111110000011111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111101110001111111111111111111111111111111111111111111111011110000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111,
160'b1110011111001111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111001111111111111111111111111111111111111111111111111000000000000000000000110000000000111111111111111111111111111111111111111111111111111111111111111111,
160'b1001111111000001001111111111111111111111111111111111111111111000000000000000000001111000000000011111111111111111111111111111111111111111111111111111111111111111,
160'b0001111111000001000011101111111111111111111111111111111111111110000000000000000011111110000000000111111111111111111111111111111111111111111111111111111111111111,
160'b0001111111000001100011100011111111111111111111111111111111111111100000000000000011110111100000000011111111111111111111111111111111111111111111111111111111111111,
160'b0000111111000001110011100001111111111111111111111111111111111111100000000111111111000111110000000001111111111111111111111111001111111111111111111111111111111111,
160'b1111001111110011111111110001111111111111111111111111111111111111100000001111111111011111100000000001111111111111111111111000000111111111111111111111111111111111,
160'b1111100111111011111111111110011111111111111111111111111111111111111111111111111111111111111011100001111111111111111111111000001111111111111111111111111111111111,
160'b1111100111110011111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111100011111111111111111111111111111111111,
160'b0111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111,
160'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111,
160'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111,
160'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111,
160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111,
160'b1111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
160'b1111111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111,
160'b1111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111,
160'b1111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111,
160'b1111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111,
160'b1111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111,
160'b1111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111,
160'b1111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000100000000011111111111111111111111,
160'b1111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111111111111110011111111100000000000000001100000111111111111111111111,
160'b1111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111000000111111100000000000000001110000011111111111111111111,
160'b1111111111111111111111111111100000000000000000000000000000011111111111111111111111111111111111111111000000000011100000000000000000001110000000111111111111111111,
160'b1111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000001111000000011111111111111111,
160'b1111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000001111000000000001111111111111111,
160'b1111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000011110011111000000100001111111111111111,
160'b1111111111111111111111111100000000000000000000000000001111111111111111111111111111001111000000000000000000000000000000100011111111111000011000111111111111111111,
160'b1111111111111111111111111000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000011110000111111110000111000111111111111111111,
160'b1111111111111111111111110000000000000000000000000000111111111111111111111111111000000000000000000000000110000000001111000001111111110011110001111111111111111111,
160'b1111111111111111111111100000000000000000000000000001111111111111111111111111110000000000000000000000001100000001111000000011111111100111100011111111111111111111,
160'b1111111111111111111111000000000000000000000000000011111111111111111111111111100000000000000000000000011100000011111000001111111111000111000111111111111111111111,
160'b1111111111111111111110000000000000000000000000000111111111111111111111111111000000000000000000000000111000000111110000011111111110001110001111111111111111111111,
160'b1111111111111111111110000000000000000000000000001111111111111111111111111111000000000000000000000001110000001111110000111111111110001111111111111111111111111111,
160'b1111111111111111111100000000000000000000000000011111111111111111111111111110001011001100000000000001100000111111110011111111111100011111111111111111111111111111,
160'b1111111111111111111100000000000000000000010000111111111111111111111111111100011111111110001100000011100011111111100011111111111100111111111111111111111111111111,
160'b1111111111111111111000000000000000000000000001111111111111111111111111111000111111111110001110000111000111111111100111111111111101111111111111111111111111111111,
160'b1111111111111111110000000000000000000001000011111111111111111111111111110001111111111110001110001111001111111111000111111111111011111111111111111111111111111111,
160'b1111111111111111110000000000000000000010000111111111111111111111111111110011111111111110001111111110011111111111011111111111111111111111111111111111111001111111,
160'b1111111111111111100000000000000000000100001111111111111111111111111111101111111111111110000111111111111111111110111111111111111111111111111111111111110011111111,
160'b1111111111111111100000000000000000000000011111111111111111111111111111001111111111111111000000011111111111111111111111101111111111111111111111111111100011111111,
160'b1111111111111111000000000000000000000000111111111111111111111111111100011111111111111111100000000111111111111111111111001111111111111111111111111111100111111111
};

reg pixel;


wire display_en;
//reg [9:0] h_count;
wire [11:0] h_count;
//reg [9:0] v_count;
wire [11:0] v_count;



localparam h_pixel_max = 800; 
localparam v_pixel_max = 600; 
localparam h_pixel_half = 400; 
localparam v_pixel_half = 300;

    
reg [4:0] addr;	
reg [7:0] data;	
reg [7:0] data_out;
always@(addr) begin
	case (addr)
		
		0 : data =  0;
		1 : data = 16;
		2 : data = 31;
		3 : data = 45;
		4 : data = 58;
 		5 : data = 67;
  		6 : data = 74;
		7 : data = 77;
		8 : data = 77;
		9 : data = 74;
		10 : data = 67;
		11 : data = 58;
		12 : data = 45;
		13 : data = 31;
		14 : data = 16;
		15 : data = 0;
		16 : data = -16;
		17 : data = -31;
		18 : data = -45;
		19 : data = -58;
		20 : data = -67;
		21 : data = -74;
		22 : data = -77;
		23 : data = -77;
  		24 : data = -74;
		25 : data = -67;
		26 : data = -58;
		27 : data = -45;
		28 : data = -31;
		29 : data = -16;
		default : data =  0;
	endcase
end

reg[22:0] div_cntr1;
reg[22:0] div_cntr2;     
reg half_sec_pulse;                  

always@(posedge clk_in)
begin
	div_cntr1 <= div_cntr1 + 1;
		if (div_cntr1 == 0)
					if (div_cntr2 == 0)
								   begin
									   div_cntr2 <= 0;
									   half_sec_pulse <= 1; 
								   end
					else
					    div_cntr2 <= div_cntr2 + 1;
		else
			half_sec_pulse <= 0;                            
		   
end    


always @(posedge half_sec_pulse) begin

        data_out <= data;
        addr <= addr + 1;
        if(addr == 29)
            addr <= 0;

end

// FOR AUDIO IN INTERACTION
assign red_led = analog_in;
assign green_led = analog_in;  

// FOR KEY INTERACTION key[8:0]

// FOR POT INTERACTION

reg [15:0] adc_count= 0; //16 bits to count how long it's taking to charge. 32,768 is the max value. 1 extra MSB bit for just discharging the cap.
reg [14:0] pot_value= 0; //to store cap charge time value
reg [14:0] final_pot_value= 0;

wire adc_in;
reg adc_sample = 1; //first time through we want to sample the cap value

wire adc;


assign pot_in = (adc_sample) ? 1'bZ : 1'b0;
assign adc_in = pot_in;

// for a 25MHz clock we divide 100MHz by 4
reg [1:0] clk_div = 0;

always @(posedge clk_in)
begin
     clk_div <= clk_div + 1;
end


always @(posedge clk_div[1]) begin //25MHz clock
	
	adc_count <= adc_count + 1; // start counting

		if(adc_count>=16'b1000000000000000 )begin // once we have rolled over 15 bit counter...

			adc_sample <= 1'b0; // ...discharge cap for a while to restart the process.

		end

		else begin
			
			adc_sample<=1'b1; //put cap pin in high 'Z'

			if(adc_in==1'b1) begin // if cap charged...

				pot_value[14:0]<=adc_count[14:0]; //store this value in pot 

				
			end

		end

end


// FOR SOUND INTERACTION 

// FOR AUDIO IN INTERACTION

//Check if we can create RGB colors
always @(posedge clk_in) begin
			
	if (display_en) begin
	
		//divide hc (once in visible area) by 8, divide vc (once in visible area) by 8 and multiply by the row width
		pixel = heart[(((h_count)>>(~key[7:4]))+(((v_count)>>(~key[3:0]))*160))];
			
				if (pixel == 1'b1) begin
				//yellow
					r_out <= key[2:0];
					g_out <= key[5:3];
					b_out <= key[8:6];	
				end
				else begin
					r_out <= key[8:6];
					g_out <= key[5:3];
					b_out <= key[2:0];
				end
	end

	else begin
	
		r_out <= 3'b000;
	    g_out <= 3'b000;
		b_out <= 3'b000;	
			
	end	

end
vga_sync vga_s(
      .clk_in(clk_div[0]),         //50MHz
      .h_sync(h_sync),
      .v_sync(v_sync),
      .h_count(h_count),
      .v_count(v_count),
      .display_en(display_en) // '1' => pixel region
      );

endmodule
